** Generated for: hspiceD
** Generated on: Sep 24 04:30:05 2023
** Design library name: yaoyuan
** Design cell name: tb_OTA_two
** Design view name: config
.GLOBAL vdd!
.PARAM cap=1.5e-12 i1=1.5e-05 i2=1.5e-05 l=5e-07 r=1000


.TEMP 25
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2
+    HIER_DELIM=0


.LIB "D:/paperwork/smic18/models/hspice/ms018_enhanced_v1p11.lib" TT
.LIB "D:/paperwork/smic18/models/hspice/ms018_enhanced_v1p11.lib" BJT_TT
.LIB "D:/paperwork/smic18/models/hspice/ms018_enhanced_v1p11.lib" DIO_TT
.LIB "D:/paperwork/smic18/models/hspice/ms018_enhanced_v1p11.lib" RES_TT
.LIB "D:/paperwork/smic18/models/hspice/ms018_enhanced_v1p11.lib" MIM_TT
.LIB "D:/paperwork/smic18/models/hspice/ms018_enhanced_v1p11.lib" VAR_TT
.LIB "D:/paperwork/smic18/models/hspice/mse018_v1p11_rf.lib" TT
.LIB "D:/paperwork/smic18/models/hspice/mse018_v1p11_rf.lib" RES_TT
.LIB "D:/paperwork/smic18/models/hspice/mse018_v1p11_rf.lib" MIM_TT
.LIB "D:/paperwork/smic18/models/hspice/mse018_v1p11_rf.lib" VAR_TT
.LIB "D:/paperwork/smic18/models/hspice/mse018_v1p11_rf.lib" IND_RF_PSUB_TT
.LIB "D:/paperwork/smic18/models/hspice/mse018_v1p11_rf.lib" IND_RF_TT
.LIB "D:/paperwork/smic18/models/hspice/mse018_v1p11_rf.lib" 3TDIFF_PSUB_TT
.LIB "D:/paperwork/smic18/models/hspice/mse018_v1p11_rf.lib" 3TDIFF_TT
.LIB "D:/paperwork/smic18/models/hspice/mse018_v1p11_rf.lib" 2TDIFF_PSUB_TT
.LIB "D:/paperwork/smic18/models/hspice/mse018_v1p11_rf.lib" 2TDIFF_TT

** Library name: yaoyuan
** Cell name: OTA_two
** View name: schematic
** Inherited view list: spectre spice verilog behavioral functional hdl system verilogNetlist schematic cmos.sch cmos_sch veriloga ahdl
.subckt OTA_two ibias1 ibias2 out _net0 _net1
mnm9 ibias2 ibias2 0 0 n18 m=1 w=13.5e-6 l=1e-6 nf=1 ad=6.48e-12 as=6.48e-12 pd=27.96e-6 ps=27.96e-6 nrd=20e-3 nrs=20e-3 sa=480e-9 sb=480e-9 sd=0 sca=0 scb=0 scc=0
mnm5 net3 _net0 net1 0 n18 m=1 w='(6uL)' l=l nf=1 ad='(((6uL) / (1)) < 419.5n) ? ((int((1) / 2.0) * (((220n + 200n) * 420n) + (((6uL) / (1)) * 200n))) + ((((1) / 2) - int((1) / 2) != 0) ? (((220n > (220n + 200n) ? 220n : (220n + 200n)) * 420n) + (((6uL) / (1)) * 100n)) : 0)) / 1 : ((int((1) / 2.0) * ((220n + 320n) * ((6uL) / (1)))) + ((((1) / 2) - int((1) / 2) != 0) ? ((320n > (220n + 260n) ? 320n : (220n + 260n)) * ((6uL) / (1))) : 0)) / 1' as='(((6uL) / (1)) < 419.5n) ? ((((220n > (220n + 200n) ? 220n : (220n + 200n)) * 420n) + (((6uL) / (1)) * 100n)) + (0 * ((((6uL) / (1)) < 419.5n) ? 420n : ((6uL) / (1)))) + (int(((1) - 1) / 2.0) * (((220n + 200n) * 420n) + (((6uL) / (1)) * 200n))) + ((((1) / 2) - int((1) / 2) == 0) ? (((220n > (220n + 200n) ? 220n : (220n + 200n)) * 420n) + (((6uL) / (1)) * 100n)) : 0)) / 1 : (((320n > (220n + 260n) ? 320n : (220n + 260n)) * ((6uL) / (1))) + (0 * ((((6uL) / (1)) < 419.5n) ? 420n : ((6uL) / (1)))) + (int(((1) - 1) / 2.0) * ((220n + 320n) * ((6uL) / (1)))) + ((((1) / 2) - 
+int((1) / 2) == 0) ? ((320n > (220n + 260n) ? 320n : (220n + 260n)) * ((6uL) / (1))) : 0)) / 1' pd='(((6uL) / (1)) < 419.5n) ? ((int((1) / 2.0) * ((2 * (220n + 200n)) + 1.24u)) + ((((1) / 2) - int((1) / 2) != 0) ? ((2 * (220n > (220n + 200n) ? 220n : (220n + 200n))) + 1.04u) : 0)) / 1 : ((int((1) / 2.0) * ((2 * (220n + 320n)) + (2 * ((6uL) / (1))))) + ((((1) / 2) - int((1) / 2) != 0) ? ((2 * (320n > (220n + 260n) ? 320n : (220n + 260n))) + (2 * ((6uL) / (1)))) : 0)) / 1' ps='(((6uL) / (1)) < 419.5n) ? (((2 * (220n > (220n + 200n) ? 220n : (220n + 200n))) + 1.04u) + 0 + (int(((1) - 1) / 2.0) * ((2 * (220n + 200n)) + 1.24u)) + ((((1) / 2) - int((1) / 2) == 0) ? ((2 * (220n > (220n + 200n) ? 220n : (220n + 200n))) + 1.04u) : 0)) / 1 : (((2 * (320n > (220n + 260n) ? 320n : (220n + 260n))) + (2 * ((6uL) / (1)))) + 0 + (int(((1) - 1) / 2.0) * ((2 * (220n + 320n)) + (2 * ((6uL) / (1))))) + ((((1) / 2) - int((1) / 2) == 0) ? ((2 * (320n > (220n + 260n) ? 320n : (220n + 260n))) + (2 * ((6uL) / (1)))) : 0)) / 1'
+nrd='( 2.2e-07/2 + 1.6e-07) / (((6uL) / (1)) * (1))' nrs='( 2.2e-07/2 + 1.6e-07) / (((6uL) / (1)) * (1))' sa='(((6uL) / (1)) < 419.5n) ? (220n > (220n + 200n) ? 220n : (220n + 200n)) + 1e-07 : (320n > (220n + 260n) ? 320n : (220n + 260n))' sb='(((6uL) / (1)) < 419.5n) ? (220n > (220n + 200n) ? 220n : (220n + 200n)) + 1e-07 : (320n > (220n + 260n) ? 320n : (220n + 260n))' sd=0 sca=0 scb=0 scc=0
mnm4 net2 _net1 net1 0 n18 m=1 w='(6uL)' l=l nf=1 ad='(((6uL) / (1)) < 419.5n) ? ((int((1) / 2.0) * (((220n + 200n) * 420n) + (((6uL) / (1)) * 200n))) + ((((1) / 2) - int((1) / 2) != 0) ? (((220n > (220n + 200n) ? 220n : (220n + 200n)) * 420n) + (((6uL) / (1)) * 100n)) : 0)) / 1 : ((int((1) / 2.0) * ((220n + 320n) * ((6uL) / (1)))) + ((((1) / 2) - int((1) / 2) != 0) ? ((320n > (220n + 260n) ? 320n : (220n + 260n)) * ((6uL) / (1))) : 0)) / 1' as='(((6uL) / (1)) < 419.5n) ? ((((220n > (220n + 200n) ? 220n : (220n + 200n)) * 420n) + (((6uL) / (1)) * 100n)) + (0 * ((((6uL) / (1)) < 419.5n) ? 420n : ((6uL) / (1)))) + (int(((1) - 1) / 2.0) * (((220n + 200n) * 420n) + (((6uL) / (1)) * 200n))) + ((((1) / 2) - int((1) / 2) == 0) ? (((220n > (220n + 200n) ? 220n : (220n + 200n)) * 420n) + (((6uL) / (1)) * 100n)) : 0)) / 1 : (((320n > (220n + 260n) ? 320n : (220n + 260n)) * ((6uL) / (1))) + (0 * ((((6uL) / (1)) < 419.5n) ? 420n : ((6uL) / (1)))) + (int(((1) - 1) / 2.0) * ((220n + 320n) * ((6uL) / (1)))) + ((((1) / 2) - 
+int((1) / 2) == 0) ? ((320n > (220n + 260n) ? 320n : (220n + 260n)) * ((6uL) / (1))) : 0)) / 1' pd='(((6uL) / (1)) < 419.5n) ? ((int((1) / 2.0) * ((2 * (220n + 200n)) + 1.24u)) + ((((1) / 2) - int((1) / 2) != 0) ? ((2 * (220n > (220n + 200n) ? 220n : (220n + 200n))) + 1.04u) : 0)) / 1 : ((int((1) / 2.0) * ((2 * (220n + 320n)) + (2 * ((6uL) / (1))))) + ((((1) / 2) - int((1) / 2) != 0) ? ((2 * (320n > (220n + 260n) ? 320n : (220n + 260n))) + (2 * ((6uL) / (1)))) : 0)) / 1' ps='(((6uL) / (1)) < 419.5n) ? (((2 * (220n > (220n + 200n) ? 220n : (220n + 200n))) + 1.04u) + 0 + (int(((1) - 1) / 2.0) * ((2 * (220n + 200n)) + 1.24u)) + ((((1) / 2) - int((1) / 2) == 0) ? ((2 * (220n > (220n + 200n) ? 220n : (220n + 200n))) + 1.04u) : 0)) / 1 : (((2 * (320n > (220n + 260n) ? 320n : (220n + 260n))) + (2 * ((6uL) / (1)))) + 0 + (int(((1) - 1) / 2.0) * ((2 * (220n + 320n)) + (2 * ((6uL) / (1))))) + ((((1) / 2) - int((1) / 2) == 0) ? ((2 * (320n > (220n + 260n) ? 320n : (220n + 260n))) + (2 * ((6uL) / (1)))) : 0)) / 1'
+nrd='( 2.2e-07/2 + 1.6e-07) / (((6uL) / (1)) * (1))' nrs='( 2.2e-07/2 + 1.6e-07) / (((6uL) / (1)) * (1))' sa='(((6uL) / (1)) < 419.5n) ? (220n > (220n + 200n) ? 220n : (220n + 200n)) + 1e-07 : (320n > (220n + 260n) ? 320n : (220n + 260n))' sb='(((6uL) / (1)) < 419.5n) ? (220n > (220n + 200n) ? 220n : (220n + 200n)) + 1e-07 : (320n > (220n + 260n) ? 320n : (220n + 260n))' sd=0 sca=0 scb=0 scc=0
mnm3 out ibias2 0 0 n18 m=1 w=81e-6 l=1e-6 nf=1 ad=38.88e-12 as=38.88e-12 pd=162.96e-6 ps=162.96e-6 nrd=3.33333e-3 nrs=3.33333e-3 sa=480e-9 sb=480e-9 sd=0 sca=0 scb=0 scc=0
mnm2 net1 ibias1 0 0 n18 m=1 w='(13.5uL)' l=l nf=1 ad='(((13.5uL) / (1)) < 419.5n) ? ((int((1) / 2.0) * (((220n + 200n) * 420n) + (((13.5uL) / (1)) * 200n))) + ((((1) / 2) - int((1) / 2) != 0) ? (((220n > (220n + 200n) ? 220n : (220n + 200n)) * 420n) + (((13.5uL) / (1)) * 100n)) : 0)) / 1 : ((int((1) / 2.0) * ((220n + 320n) * ((13.5uL) / (1)))) + ((((1) / 2) - int((1) / 2) != 0) ? ((320n > (220n + 260n) ? 320n : (220n + 260n)) * ((13.5uL) / (1))) : 0)) / 1' as='(((13.5uL) / (1)) < 419.5n) ? ((((220n > (220n + 200n) ? 220n : (220n + 200n)) * 420n) + (((13.5uL) / (1)) * 100n)) + (0 * ((((13.5uL) / (1)) < 419.5n) ? 420n : ((13.5uL) / (1)))) + (int(((1) - 1) / 2.0) * (((220n + 200n) * 420n) + (((13.5uL) / (1)) * 200n))) + ((((1) / 2) - int((1) / 2) == 0) ? (((220n > (220n + 200n) ? 220n : (220n + 200n)) * 420n) + (((13.5uL) / (1)) * 100n)) : 0)) / 1 : (((320n > (220n + 260n) ? 320n : (220n + 260n)) * ((13.5uL) / (1))) + (0 * ((((13.5uL) / (1)) < 419.5n) ? 420n : ((13.5uL) / (1)))) + (int(((1) - 1) / 2.0) *
+((220n + 320n) * ((13.5uL) / (1)))) + ((((1) / 2) - int((1) / 2) == 0) ? ((320n > (220n + 260n) ? 320n : (220n + 260n)) * ((13.5uL) / (1))) : 0)) / 1' pd='(((13.5uL) / (1)) < 419.5n) ? ((int((1) / 2.0) * ((2 * (220n + 200n)) + 1.24u)) + ((((1) / 2) - int((1) / 2) != 0) ? ((2 * (220n > (220n + 200n) ? 220n : (220n + 200n))) + 1.04u) : 0)) / 1 : ((int((1) / 2.0) * ((2 * (220n + 320n)) + (2 * ((13.5uL) / (1))))) + ((((1) / 2) - int((1) / 2) != 0) ? ((2 * (320n > (220n + 260n) ? 320n : (220n + 260n))) + (2 * ((13.5uL) / (1)))) : 0)) / 1' ps='(((13.5uL) / (1)) < 419.5n) ? (((2 * (220n > (220n + 200n) ? 220n : (220n + 200n))) + 1.04u) + 0 + (int(((1) - 1) / 2.0) * ((2 * (220n + 200n)) + 1.24u)) + ((((1) / 2) - int((1) / 2) == 0) ? ((2 * (220n > (220n + 200n) ? 220n : (220n + 200n))) + 1.04u) : 0)) / 1 : (((2 * (320n > (220n + 260n) ? 320n : (220n + 260n))) + (2 * ((13.5uL) / (1)))) + 0 + (int(((1) - 1) / 2.0) * ((2 * (220n + 320n)) + (2 * ((13.5uL) / (1))))) + ((((1) / 2) - int((1) / 2) == 0) ? ((2 * (320n >
+(220n + 260n) ? 320n : (220n + 260n))) + (2 * ((13.5uL) / (1)))) : 0)) / 1' nrd='( 2.2e-07/2 + 1.6e-07) / (((13.5uL) / (1)) * (1))' nrs='( 2.2e-07/2 + 1.6e-07) / (((13.5uL) / (1)) * (1))' sa='(((13.5uL) / (1)) < 419.5n) ? (220n > (220n + 200n) ? 220n : (220n + 200n)) + 1e-07 : (320n > (220n + 260n) ? 320n : (220n + 260n))' sb='(((13.5uL) / (1)) < 419.5n) ? (220n > (220n + 200n) ? 220n : (220n + 200n)) + 1e-07 : (320n > (220n + 260n) ? 320n : (220n + 260n))' sd=0 sca=0 scb=0 scc=0
mnm1 ibias1 ibias1 0 0 n18 m=1 w=13.5e-6 l=1e-6 nf=1 ad=6.48e-12 as=6.48e-12 pd=27.96e-6 ps=27.96e-6 nrd=20e-3 nrs=20e-3 sa=480e-9 sb=480e-9 sd=0 sca=0 scb=0 scc=0
mpm0 net2 net2 vdd! vdd! p18 m=1 w='(3.5uL)' l=l nf=1 ad='(((3.5uL) / (1)) < 419.5n) ? ((int((1) / 2.0) * (((220n + 200n) * 420n) + (((3.5uL) / (1)) * 200n))) + ((((1) / 2) - int((1) / 2) != 0) ? (((220n > (220n + 200n) ? 220n : (220n + 200n)) * 420n) + (((3.5uL) / (1)) * 100n)) : 0)) / 1 : ((int((1) / 2.0) * ((220n + 320n) * ((3.5uL) / (1)))) + ((((1) / 2) - int((1) / 2) != 0) ? ((320n > (220n + 260n) ? 320n : (220n + 260n)) * ((3.5uL) / (1))) : 0)) / 1' as='(((3.5uL) / (1)) < 419.5n) ? ((((220n > (220n + 200n) ? 220n : (220n + 200n)) * 420n) + (((3.5uL) / (1)) * 100n)) + (0 * ((((3.5uL) / (1)) < 419.5n) ? 420n : ((3.5uL) / (1)))) + (int(((1) - 1) / 2.0) * (((220n + 200n) * 420n) + (((3.5uL) / (1)) * 200n))) + ((((1) / 2) - int((1) / 2) == 0) ? (((220n > (220n + 200n) ? 220n : (220n + 200n)) * 420n) + (((3.5uL) / (1)) * 100n)) : 0)) / 1 : (((320n > (220n + 260n) ? 320n : (220n + 260n)) * ((3.5uL) / (1))) + (0 * ((((3.5uL) / (1)) < 419.5n) ? 420n : ((3.5uL) / (1)))) + (int(((1) - 1) / 2.0) * ((220n + 320n) * 
+((3.5uL) / (1)))) + ((((1) / 2) - int((1) / 2) == 0) ? ((320n > (220n + 260n) ? 320n : (220n + 260n)) * ((3.5uL) / (1))) : 0)) / 1' pd='(((3.5uL) / (1)) < 419.5n) ? ((int((1) / 2.0) * ((2 * (220n + 200n)) + 1.24u)) + ((((1) / 2) - int((1) / 2) != 0) ? ((2 * (220n > (220n + 200n) ? 220n : (220n + 200n))) + 1.04u) : 0)) / 1 : ((int((1) / 2.0) * ((2 * (220n + 320n)) + (2 * ((3.5uL) / (1))))) + ((((1) / 2) - int((1) / 2) != 0) ? ((2 * (320n > (220n + 260n) ? 320n : (220n + 260n))) + (2 * ((3.5uL) / (1)))) : 0)) / 1' ps='(((3.5uL) / (1)) < 419.5n) ? (((2 * (220n > (220n + 200n) ? 220n : (220n + 200n))) + 1.04u) + 0 + (int(((1) - 1) / 2.0) * ((2 * (220n + 200n)) + 1.24u)) + ((((1) / 2) - int((1) / 2) == 0) ? ((2 * (220n > (220n + 200n) ? 220n : (220n + 200n))) + 1.04u) : 0)) / 1 : (((2 * (320n > (220n + 260n) ? 320n : (220n + 260n))) + (2 * ((3.5uL) / (1)))) + 0 + (int(((1) - 1) / 2.0) * ((2 * (220n + 320n)) + (2 * ((3.5uL) / (1))))) + ((((1) / 2) - int((1) / 2) == 0) ? ((2 * (320n > (220n + 260n) ? 320n : (220n
++ 260n))) + (2 * ((3.5uL) / (1)))) : 0)) / 1' nrd='( 2.2e-07/2 + 1.6e-07) / (((3.5uL) / (1)) * (1))' nrs='( 2.2e-07/2 + 1.6e-07) / (((3.5uL) / (1)) * (1))' sa='(((3.5uL) / (1)) < 419.5n) ? (220n > (220n + 200n) ? 220n : (220n + 200n)) + 1e-07 : (320n > (220n + 260n) ? 320n : (220n + 260n))' sb='(((3.5uL) / (1)) < 419.5n) ? (220n > (220n + 200n) ? 220n : (220n + 200n)) + 1e-07 : (320n > (220n + 260n) ? 320n : (220n + 260n))' sd=0 sca=0 scb=0 scc=0
mpm2 out net3 vdd! vdd! p18 m=1 w=45e-6 l=1e-6 nf=1 ad=21.6e-12 as=21.6e-12 pd=90.96e-6 ps=90.96e-6 nrd=6e-3 nrs=6e-3 sa=480e-9 sb=480e-9 sd=0 sca=0 scb=0 scc=0
mpm1 net3 net2 vdd! vdd! p18 m=1 w='(3.5uL)' l=l nf=1 ad='(((3.5uL) / (1)) < 419.5n) ? ((int((1) / 2.0) * (((220n + 200n) * 420n) + (((3.5uL) / (1)) * 200n))) + ((((1) / 2) - int((1) / 2) != 0) ? (((220n > (220n + 200n) ? 220n : (220n + 200n)) * 420n) + (((3.5uL) / (1)) * 100n)) : 0)) / 1 : ((int((1) / 2.0) * ((220n + 320n) * ((3.5uL) / (1)))) + ((((1) / 2) - int((1) / 2) != 0) ? ((320n > (220n + 260n) ? 320n : (220n + 260n)) * ((3.5uL) / (1))) : 0)) / 1' as='(((3.5uL) / (1)) < 419.5n) ? ((((220n > (220n + 200n) ? 220n : (220n + 200n)) * 420n) + (((3.5uL) / (1)) * 100n)) + (0 * ((((3.5uL) / (1)) < 419.5n) ? 420n : ((3.5uL) / (1)))) + (int(((1) - 1) / 2.0) * (((220n + 200n) * 420n) + (((3.5uL) / (1)) * 200n))) + ((((1) / 2) - int((1) / 2) == 0) ? (((220n > (220n + 200n) ? 220n : (220n + 200n)) * 420n) + (((3.5uL) / (1)) * 100n)) : 0)) / 1 : (((320n > (220n + 260n) ? 320n : (220n + 260n)) * ((3.5uL) / (1))) + (0 * ((((3.5uL) / (1)) < 419.5n) ? 420n : ((3.5uL) / (1)))) + (int(((1) - 1) / 2.0) * ((220n + 320n) * 
+((3.5uL) / (1)))) + ((((1) / 2) - int((1) / 2) == 0) ? ((320n > (220n + 260n) ? 320n : (220n + 260n)) * ((3.5uL) / (1))) : 0)) / 1' pd='(((3.5uL) / (1)) < 419.5n) ? ((int((1) / 2.0) * ((2 * (220n + 200n)) + 1.24u)) + ((((1) / 2) - int((1) / 2) != 0) ? ((2 * (220n > (220n + 200n) ? 220n : (220n + 200n))) + 1.04u) : 0)) / 1 : ((int((1) / 2.0) * ((2 * (220n + 320n)) + (2 * ((3.5uL) / (1))))) + ((((1) / 2) - int((1) / 2) != 0) ? ((2 * (320n > (220n + 260n) ? 320n : (220n + 260n))) + (2 * ((3.5uL) / (1)))) : 0)) / 1' ps='(((3.5uL) / (1)) < 419.5n) ? (((2 * (220n > (220n + 200n) ? 220n : (220n + 200n))) + 1.04u) + 0 + (int(((1) - 1) / 2.0) * ((2 * (220n + 200n)) + 1.24u)) + ((((1) / 2) - int((1) / 2) == 0) ? ((2 * (220n > (220n + 200n) ? 220n : (220n + 200n))) + 1.04u) : 0)) / 1 : (((2 * (320n > (220n + 260n) ? 320n : (220n + 260n))) + (2 * ((3.5uL) / (1)))) + 0 + (int(((1) - 1) / 2.0) * ((2 * (220n + 320n)) + (2 * ((3.5uL) / (1))))) + ((((1) / 2) - int((1) / 2) == 0) ? ((2 * (320n > (220n + 260n) ? 320n : (220n
++ 260n))) + (2 * ((3.5uL) / (1)))) : 0)) / 1' nrd='( 2.2e-07/2 + 1.6e-07) / (((3.5uL) / (1)) * (1))' nrs='( 2.2e-07/2 + 1.6e-07) / (((3.5uL) / (1)) * (1))' sa='(((3.5uL) / (1)) < 419.5n) ? (220n > (220n + 200n) ? 220n : (220n + 200n)) + 1e-07 : (320n > (220n + 260n) ? 320n : (220n + 260n))' sb='(((3.5uL) / (1)) < 419.5n) ? (220n > (220n + 200n) ? 220n : (220n + 200n)) + 1e-07 : (320n > (220n + 260n) ? 320n : (220n + 260n))' sd=0 sca=0 scb=0 scc=0
c0 net3 net6 {cap}
r0 net6 out {r}
.ends OTA_two
** End of subcircuit definition.

** Library name: yaoyuan
** Cell name: tb_OTA_two
** View name: schematic
** Inherited view list: spectre spice verilog behavioral functional hdl system verilogNetlist schematic cmos.sch cmos_sch veriloga ahdl
xi0 ibias1 ibias2 net4 net2 net5 OTA_two
v4 net2 0 DC=900e-3 AC 0.5 180
v5 net5 0 DC=900e-3 AC 0.5 0
vi vdd! 0 DC=1.8
i9 vdd! ibias2 DC=i2
i3 vdd! ibias1 DC=i1
c0 net4 0 10e-12

.control 
AC DEC 10 0.01 100000K
op
.endc

.END
